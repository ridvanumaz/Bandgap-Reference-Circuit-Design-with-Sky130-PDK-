magic
tech sky130A
magscale 1 2
timestamp 1670911998
<< nwell >>
rect -13300 8300 27760 10700
<< mvnmos >>
rect -12200 3700 -11700 5700
rect -11200 3700 -10700 5700
rect -10200 3700 -9700 5700
rect -9200 3700 -8700 5700
rect -7200 3700 -7000 5700
rect -6500 3700 -6300 5700
rect -5800 3700 -5600 5700
rect -5100 3700 -4900 5700
rect -3400 3700 -2400 5700
rect -1900 3700 -900 5700
rect -400 3700 600 5700
rect 2100 3700 3100 5700
rect 3600 3700 4600 5700
rect 6100 3700 7100 5700
rect 7600 3700 8600 5700
rect 10100 3700 11100 5700
rect 11600 3700 12600 5700
rect 13100 3700 14100 5700
<< mvpmos >>
rect -12200 8500 -11200 10500
rect -9700 8500 -8700 10500
rect -8200 8500 -7200 10500
rect -5700 8500 -4700 10500
rect -4200 8500 -3200 10500
rect -1700 8500 -700 10500
rect -200 8500 800 10500
rect 2300 8500 3300 10500
rect 3800 8500 4800 10500
rect 5300 8500 6300 10500
rect 7800 8500 8800 10500
rect 9300 8500 10300 10500
rect 11800 8500 12800 10500
rect 13300 8500 14300 10500
rect 15800 8500 16800 10500
rect 17300 8500 18300 10500
rect 19800 8500 20800 10500
rect 21300 8500 22300 10500
rect 22800 8500 23800 10500
rect 25300 8500 26300 10500
<< mvndiff >>
rect -12700 5520 -12200 5700
rect -12700 3840 -12540 5520
rect -12360 3840 -12200 5520
rect -12700 3700 -12200 3840
rect -11700 5520 -11200 5700
rect -11700 3840 -11540 5520
rect -11360 3840 -11200 5520
rect -11700 3700 -11200 3840
rect -10700 5520 -10200 5700
rect -10700 3840 -10540 5520
rect -10360 3840 -10200 5520
rect -10700 3700 -10200 3840
rect -9700 5520 -9200 5700
rect -9700 3840 -9540 5520
rect -9360 3840 -9200 5520
rect -9700 3700 -9200 3840
rect -8700 5520 -8200 5700
rect -8700 3840 -8540 5520
rect -8360 3840 -8200 5520
rect -7700 5520 -7200 5700
rect -8700 3700 -8200 3840
rect -7700 3840 -7540 5520
rect -7360 3840 -7200 5520
rect -7700 3700 -7200 3840
rect -7000 5520 -6500 5700
rect -7000 3840 -6840 5520
rect -6660 3840 -6500 5520
rect -7000 3700 -6500 3840
rect -6300 5520 -5800 5700
rect -6300 3840 -6140 5520
rect -5960 3840 -5800 5520
rect -6300 3700 -5800 3840
rect -5600 5520 -5100 5700
rect -5600 3840 -5440 5520
rect -5260 3840 -5100 5520
rect -5600 3700 -5100 3840
rect -4900 5520 -4400 5700
rect -4900 3840 -4740 5520
rect -4560 3840 -4400 5520
rect -3900 5520 -3400 5700
rect -4900 3700 -4400 3840
rect -3900 3840 -3740 5520
rect -3560 3840 -3400 5520
rect -3900 3700 -3400 3840
rect -2400 5520 -1900 5700
rect -2400 3840 -2240 5520
rect -2060 3840 -1900 5520
rect -2400 3700 -1900 3840
rect -900 5520 -400 5700
rect -900 3840 -740 5520
rect -560 3840 -400 5520
rect -900 3700 -400 3840
rect 600 5520 1100 5700
rect 600 3840 760 5520
rect 940 3840 1100 5520
rect 1600 5520 2100 5700
rect 600 3700 1100 3840
rect 1600 3840 1760 5520
rect 1940 3840 2100 5520
rect 1600 3700 2100 3840
rect 3100 5520 3600 5700
rect 3100 3840 3260 5520
rect 3440 3840 3600 5520
rect 3100 3700 3600 3840
rect 4600 5520 5100 5700
rect 4600 3840 4760 5520
rect 4940 3840 5100 5520
rect 5600 5520 6100 5700
rect 4600 3700 5100 3840
rect 5600 3840 5760 5520
rect 5940 3840 6100 5520
rect 5600 3700 6100 3840
rect 7100 5520 7600 5700
rect 7100 3840 7260 5520
rect 7440 3840 7600 5520
rect 7100 3700 7600 3840
rect 8600 5520 9100 5700
rect 8600 3840 8760 5520
rect 8940 3840 9100 5520
rect 9600 5520 10100 5700
rect 8600 3700 9100 3840
rect 9600 3840 9760 5520
rect 9940 3840 10100 5520
rect 9600 3700 10100 3840
rect 11100 5520 11600 5700
rect 11100 3840 11260 5520
rect 11440 3840 11600 5520
rect 11100 3700 11600 3840
rect 12600 5520 13100 5700
rect 12600 3840 12760 5520
rect 12940 3840 13100 5520
rect 12600 3700 13100 3840
rect 14100 5520 14600 5700
rect 14100 3840 14260 5520
rect 14440 3840 14600 5520
rect 14100 3700 14600 3840
<< mvpdiff >>
rect -12700 10340 -12200 10500
rect -12700 8660 -12540 10340
rect -12360 8660 -12200 10340
rect -12700 8500 -12200 8660
rect -11200 10340 -10700 10500
rect -10200 10340 -9700 10500
rect -11200 8660 -11040 10340
rect -10860 8660 -10700 10340
rect -10200 8660 -10040 10340
rect -9860 8660 -9700 10340
rect -11200 8500 -10700 8660
rect -10200 8500 -9700 8660
rect -8700 10340 -8200 10500
rect -8700 8660 -8540 10340
rect -8360 8660 -8200 10340
rect -8700 8500 -8200 8660
rect -7200 10340 -6700 10500
rect -6200 10340 -5700 10500
rect -7200 8660 -7040 10340
rect -6860 8660 -6700 10340
rect -6200 8660 -6040 10340
rect -5860 8660 -5700 10340
rect -7200 8500 -6700 8660
rect -6200 8500 -5700 8660
rect -4700 10340 -4200 10500
rect -4700 8660 -4540 10340
rect -4360 8660 -4200 10340
rect -4700 8500 -4200 8660
rect -3200 10340 -2700 10500
rect -2200 10340 -1700 10500
rect -3200 8660 -3040 10340
rect -2860 8660 -2700 10340
rect -2200 8660 -2040 10340
rect -1860 8660 -1700 10340
rect -3200 8500 -2700 8660
rect -2200 8500 -1700 8660
rect -700 10340 -200 10500
rect -700 8660 -540 10340
rect -360 8660 -200 10340
rect -700 8500 -200 8660
rect 800 10340 1300 10500
rect 1800 10340 2300 10500
rect 800 8660 960 10340
rect 1140 8660 1300 10340
rect 1800 8660 1960 10340
rect 2140 8660 2300 10340
rect 800 8500 1300 8660
rect 1800 8500 2300 8660
rect 3300 10340 3800 10500
rect 3300 8660 3460 10340
rect 3640 8660 3800 10340
rect 3300 8500 3800 8660
rect 4800 10340 5300 10500
rect 4800 8660 4960 10340
rect 5140 8660 5300 10340
rect 4800 8500 5300 8660
rect 6300 10340 6800 10500
rect 7300 10340 7800 10500
rect 6300 8660 6460 10340
rect 6640 8660 6800 10340
rect 7300 8660 7460 10340
rect 7640 8660 7800 10340
rect 6300 8500 6800 8660
rect 7300 8500 7800 8660
rect 8800 10340 9300 10500
rect 8800 8660 8960 10340
rect 9140 8660 9300 10340
rect 8800 8500 9300 8660
rect 10300 10340 10800 10500
rect 11300 10340 11800 10500
rect 10300 8660 10460 10340
rect 10640 8660 10800 10340
rect 11300 8660 11460 10340
rect 11640 8660 11800 10340
rect 10300 8500 10800 8660
rect 11300 8500 11800 8660
rect 12800 10340 13300 10500
rect 12800 8660 12960 10340
rect 13140 8660 13300 10340
rect 12800 8500 13300 8660
rect 14300 10340 14800 10500
rect 15300 10340 15800 10500
rect 14300 8660 14460 10340
rect 14640 8660 14800 10340
rect 15300 8660 15460 10340
rect 15640 8660 15800 10340
rect 14300 8500 14800 8660
rect 15300 8500 15800 8660
rect 16800 10340 17300 10500
rect 16800 8660 16960 10340
rect 17140 8660 17300 10340
rect 16800 8500 17300 8660
rect 18300 10340 18800 10500
rect 19300 10340 19800 10500
rect 18300 8660 18460 10340
rect 18640 8660 18800 10340
rect 19300 8660 19460 10340
rect 19640 8660 19800 10340
rect 18300 8500 18800 8660
rect 19300 8500 19800 8660
rect 20800 10340 21300 10500
rect 20800 8660 20960 10340
rect 21140 8660 21300 10340
rect 20800 8500 21300 8660
rect 22300 10340 22800 10500
rect 22300 8660 22460 10340
rect 22640 8660 22800 10340
rect 22300 8500 22800 8660
rect 23800 10340 24300 10500
rect 24800 10340 25300 10500
rect 23800 8660 23960 10340
rect 24140 8660 24300 10340
rect 24800 8660 24960 10340
rect 25140 8660 25300 10340
rect 23800 8500 24300 8660
rect 24800 8500 25300 8660
rect 26300 10340 26800 10500
rect 26300 8660 26460 10340
rect 26640 8660 26800 10340
rect 26300 8500 26800 8660
<< mvndiffc >>
rect -12540 3840 -12360 5520
rect -11540 3840 -11360 5520
rect -10540 3840 -10360 5520
rect -9540 3840 -9360 5520
rect -8540 3840 -8360 5520
rect -7540 3840 -7360 5520
rect -6840 3840 -6660 5520
rect -6140 3840 -5960 5520
rect -5440 3840 -5260 5520
rect -4740 3840 -4560 5520
rect -3740 3840 -3560 5520
rect -2240 3840 -2060 5520
rect -740 3840 -560 5520
rect 760 3840 940 5520
rect 1760 3840 1940 5520
rect 3260 3840 3440 5520
rect 4760 3840 4940 5520
rect 5760 3840 5940 5520
rect 7260 3840 7440 5520
rect 8760 3840 8940 5520
rect 9760 3840 9940 5520
rect 11260 3840 11440 5520
rect 12760 3840 12940 5520
rect 14260 3840 14440 5520
<< mvpdiffc >>
rect -12540 8660 -12360 10340
rect -11040 8660 -10860 10340
rect -10040 8660 -9860 10340
rect -8540 8660 -8360 10340
rect -7040 8660 -6860 10340
rect -6040 8660 -5860 10340
rect -4540 8660 -4360 10340
rect -3040 8660 -2860 10340
rect -2040 8660 -1860 10340
rect -540 8660 -360 10340
rect 960 8660 1140 10340
rect 1960 8660 2140 10340
rect 3460 8660 3640 10340
rect 4960 8660 5140 10340
rect 6460 8660 6640 10340
rect 7460 8660 7640 10340
rect 8960 8660 9140 10340
rect 10460 8660 10640 10340
rect 11460 8660 11640 10340
rect 12960 8660 13140 10340
rect 14460 8660 14640 10340
rect 15460 8660 15640 10340
rect 16960 8660 17140 10340
rect 18460 8660 18640 10340
rect 19460 8660 19640 10340
rect 20960 8660 21140 10340
rect 22460 8660 22640 10340
rect 23960 8660 24140 10340
rect 24960 8660 25140 10340
rect 26460 8660 26640 10340
<< mvpsubdiff >>
rect -13200 5540 -12700 5700
rect -13200 3860 -13040 5540
rect -12860 3860 -12700 5540
rect -13200 3700 -12700 3860
rect -8200 5540 -7700 5700
rect -8200 3860 -8040 5540
rect -7860 3860 -7700 5540
rect -8200 3700 -7700 3860
rect -4400 5540 -3900 5700
rect -4400 3860 -4240 5540
rect -4060 3860 -3900 5540
rect -4400 3700 -3900 3860
rect 1100 5540 1600 5700
rect 1100 3860 1260 5540
rect 1440 3860 1600 5540
rect 1100 3700 1600 3860
rect 5100 5540 5600 5700
rect 5100 3860 5260 5540
rect 5440 3860 5600 5540
rect 5100 3700 5600 3860
rect 9100 5540 9600 5700
rect 9100 3860 9260 5540
rect 9440 3860 9600 5540
rect 9100 3700 9600 3860
rect 14600 5540 15100 5700
rect 14600 3860 14760 5540
rect 14940 3860 15100 5540
rect 14600 3700 15100 3860
<< mvnsubdiff >>
rect -13200 10340 -12700 10500
rect -13200 8660 -13040 10340
rect -12860 8660 -12700 10340
rect -13200 8500 -12700 8660
rect -10700 10340 -10200 10500
rect -10700 8660 -10540 10340
rect -10360 8660 -10200 10340
rect -10700 8500 -10200 8660
rect -6700 10340 -6200 10500
rect -6700 8660 -6540 10340
rect -6360 8660 -6200 10340
rect -6700 8500 -6200 8660
rect -2700 10340 -2200 10500
rect -2700 8660 -2540 10340
rect -2360 8660 -2200 10340
rect -2700 8500 -2200 8660
rect 1300 10340 1800 10500
rect 1300 8660 1460 10340
rect 1640 8660 1800 10340
rect 1300 8500 1800 8660
rect 6800 10340 7300 10500
rect 6800 8660 6960 10340
rect 7140 8660 7300 10340
rect 6800 8500 7300 8660
rect 10800 10340 11300 10500
rect 10800 8660 10960 10340
rect 11140 8660 11300 10340
rect 10800 8500 11300 8660
rect 14800 10340 15300 10500
rect 14800 8660 14960 10340
rect 15140 8660 15300 10340
rect 14800 8500 15300 8660
rect 18800 10340 19300 10500
rect 18800 8660 18960 10340
rect 19140 8660 19300 10340
rect 18800 8500 19300 8660
rect 24300 10340 24800 10500
rect 24300 8660 24460 10340
rect 24640 8660 24800 10340
rect 24300 8500 24800 8660
rect 26800 10340 27300 10500
rect 26800 8660 26960 10340
rect 27140 8660 27300 10340
rect 26800 8500 27300 8660
<< mvpsubdiffcont >>
rect -13040 3860 -12860 5540
rect -8040 3860 -7860 5540
rect -4240 3860 -4060 5540
rect 1260 3860 1440 5540
rect 5260 3860 5440 5540
rect 9260 3860 9440 5540
rect 14760 3860 14940 5540
<< mvnsubdiffcont >>
rect -13040 8660 -12860 10340
rect -10540 8660 -10360 10340
rect -6540 8660 -6360 10340
rect -2540 8660 -2360 10340
rect 1460 8660 1640 10340
rect 6960 8660 7140 10340
rect 10960 8660 11140 10340
rect 14960 8660 15140 10340
rect 18960 8660 19140 10340
rect 24460 8660 24640 10340
rect 26960 8660 27140 10340
<< poly >>
rect -12200 10500 -11200 10600
rect -9700 10500 -8700 10600
rect -8200 10500 -7200 10600
rect -5700 10500 -4700 10600
rect -4200 10500 -3200 10600
rect -1700 10500 -700 10600
rect -200 10500 800 10600
rect 2300 10500 3300 10600
rect 3800 10500 4800 10600
rect 5300 10500 6300 10600
rect 7800 10500 8800 10600
rect 9300 10500 10300 10600
rect 11800 10500 12800 10600
rect 13300 10500 14300 10600
rect 15800 10500 16800 10600
rect 17300 10500 18300 10600
rect 19800 10500 20800 10600
rect 21300 10500 22300 10600
rect 22800 10500 23800 10600
rect 25300 10500 26300 10600
rect -12200 8260 -11200 8500
rect -9700 8300 -8700 8500
rect -12200 8140 -12160 8260
rect -12040 8140 -11200 8260
rect -12200 8100 -11200 8140
rect -10200 8200 -8700 8300
rect -8200 8200 -7200 8500
rect -5700 8200 -4700 8500
rect -4200 8200 -3200 8500
rect -3100 8340 -2800 8400
rect -3100 8200 -3040 8340
rect -10200 8160 -3040 8200
rect -2860 8200 -2800 8340
rect -2100 8340 -1800 8400
rect -2100 8200 -2040 8340
rect -2860 8160 -2040 8200
rect -1860 8200 -1800 8340
rect -1700 8200 -700 8500
rect -200 8200 800 8500
rect 2300 8200 3300 8500
rect 3800 8200 4800 8500
rect -1860 8160 4800 8200
rect -10200 8100 4800 8160
rect 5300 8200 6300 8500
rect 6900 8340 7200 8400
rect 6900 8200 6960 8340
rect 5300 8160 6960 8200
rect 7140 8200 7200 8340
rect 7800 8200 8800 8500
rect 7140 8160 8800 8200
rect 5300 8100 8800 8160
rect 9300 8360 10300 8500
rect 9300 8160 9360 8360
rect 9540 8200 10300 8360
rect 11800 8200 12800 8500
rect 13300 8200 14300 8500
rect 15800 8440 16800 8500
rect 15800 8360 16640 8440
rect 16760 8360 16800 8440
rect 15800 8200 16800 8360
rect 9540 8160 16800 8200
rect 9300 8100 16800 8160
rect 17300 8200 18300 8500
rect 18900 8340 19200 8400
rect 18900 8200 18960 8340
rect 17300 8160 18960 8200
rect 19140 8200 19200 8340
rect 19800 8200 20800 8500
rect 19140 8160 20800 8200
rect 17300 8100 20800 8160
rect 21300 8100 22300 8500
rect 22800 8100 23800 8500
rect 25300 8260 26300 8500
rect 25300 8140 26140 8260
rect 26260 8140 26300 8260
rect 25300 8100 26300 8140
rect -10200 6200 -9700 8100
rect -6240 7400 -6060 8100
rect 15800 8000 16800 8100
rect 21300 8000 23800 8100
rect 15800 7900 23800 8000
rect -6300 7340 -6000 7400
rect -6300 7160 -6240 7340
rect -6060 7160 -6000 7340
rect -6300 7100 -6000 7160
rect -12200 6060 -11700 6100
rect -12200 5940 -12160 6060
rect -12040 5940 -11700 6060
rect -12200 5700 -11700 5940
rect -11200 6000 -9700 6200
rect -6500 6540 12600 6600
rect -6500 6360 -2240 6540
rect -2080 6360 12600 6540
rect -6500 6300 12600 6360
rect -11200 5700 -10700 6000
rect -10200 5700 -9700 6000
rect -9200 6040 -7000 6100
rect -9200 6000 -8040 6040
rect -9200 5700 -8700 6000
rect -8100 5860 -8040 6000
rect -7860 6000 -7000 6040
rect -7860 5860 -7800 6000
rect -8100 5800 -7800 5860
rect -7200 5700 -7000 6000
rect -6500 5700 -6300 6300
rect -5800 5700 -5600 6300
rect -5100 6040 -2400 6100
rect -5100 6000 -4240 6040
rect -5100 5700 -4900 6000
rect -4300 5860 -4240 6000
rect -4060 6000 -2400 6040
rect -4060 5860 -4000 6000
rect -4300 5800 -4000 5860
rect -3400 5700 -2400 6000
rect -1900 5700 -900 6300
rect -400 6040 3100 6100
rect -400 6000 1260 6040
rect -400 5700 600 6000
rect 1200 5860 1260 6000
rect 1440 6000 3100 6040
rect 1440 5860 1500 6000
rect 1200 5800 1500 5860
rect 2100 5700 3100 6000
rect 3600 5700 4600 6300
rect 6100 5700 7100 6300
rect 7600 6040 11100 6100
rect 7600 6000 9260 6040
rect 7600 5700 8600 6000
rect 9200 5860 9260 6000
rect 9440 6000 11100 6040
rect 9440 5860 9500 6000
rect 9200 5800 9500 5860
rect 10100 5700 11100 6000
rect 11600 6040 12600 6300
rect 11600 5860 12360 6040
rect 12540 5860 12600 6040
rect 11600 5700 12600 5860
rect 13100 6040 14100 6100
rect 13100 5860 13860 6040
rect 14040 5860 14100 6040
rect 13100 5700 14100 5860
rect -12200 3440 -11700 3700
rect -11200 3440 -10700 3700
rect -10200 3440 -9700 3700
rect -9200 3440 -8700 3700
rect -7200 3440 -7000 3700
rect -6500 3440 -6300 3700
rect -5800 3440 -5600 3700
rect -5100 3440 -4900 3700
rect -3400 3440 -2400 3700
rect -1900 3440 -900 3700
rect -400 3440 600 3700
rect 2100 3440 3100 3700
rect 3600 3440 4600 3700
rect 6100 3440 7100 3700
rect 7600 3440 8600 3700
rect 10100 3440 11100 3700
rect 11600 3440 12600 3700
rect 13100 3440 14100 3700
<< polycont >>
rect -12160 8140 -12040 8260
rect -3040 8160 -2860 8340
rect -2040 8160 -1860 8340
rect 6960 8160 7140 8340
rect 9360 8160 9540 8360
rect 16640 8360 16760 8440
rect 18960 8160 19140 8340
rect 26140 8140 26260 8260
rect -6240 7160 -6060 7340
rect -12160 5940 -12040 6060
rect -2240 6360 -2080 6540
rect -8040 5860 -7860 6040
rect -4240 5860 -4060 6040
rect 1260 5860 1440 6040
rect 9260 5860 9440 6040
rect 12360 5860 12540 6040
rect 13860 5860 14040 6040
<< xpolycontact >>
rect 15441 5919 15511 6409
rect 15441 4379 15511 4869
rect 15761 5919 15831 6409
rect 15761 4379 15831 4869
rect 16081 5919 16151 6409
rect 16081 4379 16151 4869
rect 16401 5919 16471 6409
rect 16401 4379 16471 4869
rect 16721 5919 16791 6409
rect 16721 4379 16791 4869
rect 17041 5919 17111 6409
rect 17041 4379 17111 4869
rect 17361 5919 17431 6409
rect 17361 4379 17431 4869
rect 17681 5919 17751 6409
rect 17681 4379 17751 4869
rect 18001 5919 18071 6400
rect 18001 4379 18071 4869
rect 18321 5919 18391 6409
rect 18321 4379 18391 4869
rect 18641 5919 18711 6409
rect 18641 4379 18711 4869
rect 18961 5919 19031 6409
rect 18961 4379 19031 4869
rect 19281 5919 19351 6409
rect 19281 4379 19351 4869
rect 19601 5719 19671 6209
rect 19601 4379 19671 4869
rect 19921 5919 19991 6409
rect 19921 4379 19991 4869
rect 20241 5919 20311 6409
rect 20241 4379 20311 4869
rect 20561 5919 20631 6409
rect 20561 4379 20631 4869
<< xpolyres >>
rect 15441 4869 15511 5919
rect 15761 4869 15831 5919
rect 16081 4869 16151 5919
rect 16401 4869 16471 5919
rect 16721 4869 16791 5919
rect 17041 4869 17111 5919
rect 17361 4869 17431 5919
rect 17681 4869 17751 5919
rect 18001 4869 18071 5919
rect 18321 4869 18391 5919
rect 18641 4869 18711 5919
rect 18961 4869 19031 5919
rect 19281 4869 19351 5919
rect 19601 4869 19671 5719
rect 19921 4869 19991 5919
rect 20241 4869 20311 5919
rect 20561 4869 20631 5919
<< locali >>
rect -13100 10398 -12800 10400
rect -12600 10398 -12300 10400
rect -13102 10348 -12300 10398
rect -13102 8663 -13046 10348
rect -12860 8663 -12548 10348
rect -12362 10340 -12300 10348
rect -13102 8660 -13040 8663
rect -12860 8660 -12540 8663
rect -12360 8660 -12300 10340
rect -13102 8600 -12300 8660
rect -11100 10353 -9800 10400
rect -11100 10343 -10541 10353
rect -11100 10340 -11039 10343
rect -11100 8660 -11040 10340
rect -10853 8668 -10541 10343
rect -10355 8668 -10047 10353
rect -9861 10340 -9800 10353
rect -10853 8660 -10540 8668
rect -10360 8660 -10040 8668
rect -9860 8660 -9800 10340
rect -11100 8658 -11039 8660
rect -10853 8658 -9800 8660
rect -11100 8600 -9800 8658
rect -8600 10340 -8300 10400
rect -8600 8660 -8540 10340
rect -8360 8660 -8300 10340
rect -8600 8600 -8300 8660
rect -7100 10340 -6800 10400
rect -7100 8660 -7040 10340
rect -6860 8660 -6800 10340
rect -12540 8260 -12360 8600
rect -7100 8400 -6800 8660
rect -6600 10348 -6300 10400
rect -6600 8663 -6551 10348
rect -6365 10340 -6300 10348
rect -6600 8660 -6540 8663
rect -6360 8660 -6300 10340
rect -6600 8600 -6300 8660
rect -6100 10340 -5800 10400
rect -6100 8660 -6040 10340
rect -5860 8660 -5800 10340
rect -6100 8400 -5800 8660
rect -4600 10340 -4300 10400
rect -4600 8660 -4540 10340
rect -4360 8660 -4300 10340
rect -4600 8600 -4300 8660
rect -3100 10340 -2800 10400
rect -3100 8660 -3040 10340
rect -2860 8660 -2800 10340
rect -3100 8600 -2800 8660
rect -2600 10353 -2300 10400
rect -2600 8668 -2542 10353
rect -2356 8668 -2300 10353
rect -2600 8660 -2540 8668
rect -2360 8660 -2300 8668
rect -2600 8600 -2300 8660
rect -2100 10340 -1800 10400
rect -2100 8660 -2040 10340
rect -1860 8660 -1800 10340
rect -2100 8600 -1800 8660
rect -600 10340 -300 10400
rect -600 8660 -540 10340
rect -360 8660 -300 10340
rect -600 8600 -300 8660
rect 900 10340 1200 10400
rect 900 8660 960 10340
rect 1140 8660 1200 10340
rect -3040 8400 -2860 8600
rect -2040 8400 -1860 8600
rect 900 8400 1200 8660
rect 1400 10348 1700 10400
rect 1400 8663 1458 10348
rect 1644 8663 1700 10348
rect 1400 8660 1460 8663
rect 1640 8660 1700 8663
rect 1400 8600 1700 8660
rect 1900 10340 2200 10400
rect 1900 8660 1960 10340
rect 2140 8660 2200 10340
rect 1900 8400 2200 8660
rect 3400 10340 3700 10400
rect 3400 8660 3460 10340
rect 3640 8660 3700 10340
rect 3400 8600 3700 8660
rect 4900 10353 5200 10400
rect 4900 8668 4959 10353
rect 5145 8668 5200 10353
rect 4900 8660 4960 8668
rect 5140 8660 5200 8668
rect 4900 8600 5200 8660
rect 6400 10353 7700 10400
rect 6400 10343 6957 10353
rect 6400 8658 6454 10343
rect 6640 8668 6957 10343
rect 7143 10348 7700 10353
rect 7143 8668 7460 10348
rect 6640 8660 6960 8668
rect 7140 8660 7460 8668
rect 7646 8663 7700 10348
rect 7640 8660 7700 8663
rect 6640 8658 7700 8660
rect 6400 8600 7700 8658
rect 8900 10340 9200 10400
rect 8900 8660 8960 10340
rect 9140 8660 9200 10340
rect 8900 8600 9200 8660
rect 10400 10353 11700 10400
rect 10400 10343 11459 10353
rect 10400 8658 10458 10343
rect 10644 10340 10961 10343
rect 10644 8660 10960 10340
rect 11147 8668 11459 10343
rect 11645 8668 11700 10353
rect 11147 8660 11460 8668
rect 11640 8660 11700 8668
rect 10644 8658 10961 8660
rect 11147 8658 11700 8660
rect 10400 8600 11700 8658
rect 12900 10340 13200 10400
rect 12900 8660 12960 10340
rect 13140 8660 13200 10340
rect 12900 8600 13200 8660
rect 14400 10353 15700 10400
rect 14400 8668 14453 10353
rect 14639 10340 14956 10353
rect 15142 10348 15700 10353
rect 14640 8668 14956 10340
rect 15142 8668 15459 10348
rect 14400 8660 14460 8668
rect 14640 8660 14960 8668
rect 15140 8663 15459 8668
rect 15645 8663 15700 10348
rect 15140 8660 15460 8663
rect 15640 8660 15700 8663
rect 14400 8600 15700 8660
rect 16900 10340 17200 10400
rect 16900 8660 16960 10340
rect 17140 8660 17200 10340
rect 6960 8400 7140 8600
rect -7100 8300 -5800 8400
rect -3100 8340 -2800 8400
rect -12200 8260 -12000 8300
rect -12540 8140 -12160 8260
rect -12040 8140 -12000 8260
rect -12200 8100 -12000 8140
rect -3100 8160 -3040 8340
rect -2860 8160 -2800 8340
rect -3100 8100 -2800 8160
rect -2100 8340 -1800 8400
rect -2100 8160 -2040 8340
rect -1860 8160 -1800 8340
rect 900 8300 2200 8400
rect 6900 8340 7200 8400
rect -2100 8100 -1800 8160
rect 6900 8160 6960 8340
rect 7140 8160 7200 8340
rect 6900 8100 7200 8160
rect 8960 8360 9140 8600
rect 9300 8360 9600 8400
rect 8960 8160 9360 8360
rect 9540 8160 9600 8360
rect 8960 7900 9120 8160
rect 9300 8100 9600 8160
rect 12960 8020 13140 8600
rect 16600 8440 16800 8500
rect 16900 8440 17200 8660
rect 18400 10348 19700 10400
rect 18400 10343 18951 10348
rect 18400 8658 18457 10343
rect 18643 8663 18951 10343
rect 19137 10340 19463 10348
rect 18643 8660 18960 8663
rect 19140 8660 19460 10340
rect 19649 8663 19700 10348
rect 19640 8660 19700 8663
rect 18643 8658 19700 8660
rect 18400 8600 19700 8658
rect 20900 10348 21200 10400
rect 20900 8663 20958 10348
rect 21144 8663 21200 10348
rect 20900 8660 20960 8663
rect 21140 8660 21200 8663
rect 20900 8600 21200 8660
rect 22400 10340 22700 10400
rect 22400 8660 22460 10340
rect 22640 8660 22700 10340
rect 16600 8360 16640 8440
rect 16760 8360 17200 8440
rect 18960 8400 19140 8600
rect 16600 8300 16800 8360
rect 18900 8340 19200 8400
rect 18900 8160 18960 8340
rect 19140 8160 19200 8340
rect 18900 8100 19200 8160
rect -11560 7700 9120 7900
rect 12760 7860 13140 8020
rect -11560 6200 -11360 7700
rect -9540 6200 -9360 7700
rect 3960 7460 4260 7502
rect -740 7442 4260 7460
rect -6300 7340 -6000 7400
rect -6300 7304 -6240 7340
rect -6840 7160 -6240 7304
rect -6060 7304 -6000 7340
rect -6060 7300 -5262 7304
rect -6060 7160 -5260 7300
rect -6840 7100 -5260 7160
rect -6841 6535 -6659 7100
rect -12200 6060 -12000 6100
rect -12540 5940 -12160 6060
rect -12040 5940 -12000 6060
rect -12540 5600 -12360 5940
rect -12200 5900 -12000 5940
rect -11560 5600 -11363 6200
rect -9541 5600 -9355 6200
rect -8100 6040 -7800 6100
rect -8100 5860 -8040 6040
rect -7860 5860 -7800 6040
rect -8100 5800 -7800 5860
rect -8040 5600 -7860 5800
rect -6840 5600 -6659 6535
rect -5444 5600 -5260 7100
rect -740 7260 4020 7442
rect -2300 6540 -2000 6600
rect -2300 6360 -2240 6540
rect -2080 6360 -2000 6540
rect -2300 6300 -2000 6360
rect -4300 6040 -4000 6100
rect -4300 5860 -4240 6040
rect -4060 5860 -4000 6040
rect -4300 5800 -4000 5860
rect -4240 5600 -4060 5800
rect -2240 5600 -2060 6300
rect -740 5600 -560 7260
rect 3960 7242 4020 7260
rect 4200 7242 4260 7442
rect 3960 7202 4260 7242
rect 3960 6960 4260 7020
rect 3260 6760 4020 6960
rect 4200 6760 4260 6960
rect 1200 6040 1500 6100
rect 1200 5860 1260 6040
rect 1440 5860 1500 6040
rect 1200 5800 1500 5860
rect 1240 5600 1440 5800
rect 3260 5600 3440 6760
rect 3960 6720 4260 6760
rect 4760 5600 4940 7700
rect 5760 5600 5940 7700
rect 6600 7460 6900 7500
rect 11660 7460 11960 7502
rect 6600 7442 11960 7460
rect 6600 7440 11720 7442
rect 6600 7240 6660 7440
rect 6840 7260 11720 7440
rect 6840 7240 6900 7260
rect 6600 7200 6900 7240
rect 6600 6960 6900 7000
rect 10660 6960 10960 7002
rect 6600 6942 10960 6960
rect 6600 6940 10720 6942
rect 6600 6740 6660 6940
rect 6840 6760 10720 6940
rect 6840 6740 6900 6760
rect 6600 6700 6900 6740
rect 7260 5600 7440 6760
rect 10660 6742 10720 6760
rect 10900 6742 10960 6942
rect 10660 6702 10960 6742
rect 9200 6040 9500 6100
rect 9200 5860 9260 6040
rect 9440 5860 9500 6040
rect 9200 5800 9500 5860
rect 9240 5600 9440 5800
rect 11260 5600 11440 7260
rect 11660 7242 11720 7260
rect 11900 7242 11960 7442
rect 11660 7202 11960 7242
rect 12300 6040 12600 6100
rect 12760 6040 12940 7860
rect 15760 7800 16120 7860
rect 22400 7800 22700 8660
rect 23900 10353 25200 10400
rect 23900 10348 24459 10353
rect 23900 8663 23956 10348
rect 24142 8668 24459 10348
rect 24645 8668 24957 10353
rect 25143 8668 25200 10353
rect 24142 8663 24460 8668
rect 23900 8660 23960 8663
rect 24140 8660 24460 8663
rect 24640 8660 24960 8668
rect 25140 8660 25200 8668
rect 23900 8600 25200 8660
rect 26400 10348 27200 10400
rect 26400 8663 26452 10348
rect 26638 10343 27200 10348
rect 26638 10340 26955 10343
rect 26400 8660 26460 8663
rect 26640 8660 26955 10340
rect 26400 8658 26955 8660
rect 27141 8658 27200 10343
rect 26400 8600 27200 8658
rect 26100 8260 26300 8300
rect 26460 8260 26640 8600
rect 26100 8140 26140 8260
rect 26260 8140 26640 8260
rect 26100 8100 26300 8140
rect 15760 7780 27760 7800
rect 15760 7620 15820 7780
rect 16060 7620 27760 7780
rect 15760 7600 27760 7620
rect 15760 7540 16120 7600
rect 22400 7580 27760 7600
rect 13380 7460 13680 7500
rect 21500 7460 22100 7500
rect 13380 7440 22100 7460
rect 13380 7240 13440 7440
rect 13620 7260 21560 7440
rect 13620 7240 13680 7260
rect 13380 7200 13680 7240
rect 21500 7240 21560 7260
rect 22040 7240 22100 7440
rect 21500 7200 22100 7240
rect 22400 7140 22700 7580
rect 13380 6960 13680 7000
rect 13380 6940 18100 6960
rect 19920 6940 22700 7140
rect 13380 6740 13440 6940
rect 13620 6760 18100 6940
rect 13620 6740 13680 6760
rect 13380 6700 13680 6740
rect 15760 6600 16120 6680
rect 15760 6540 15820 6600
rect 16060 6540 16120 6600
rect 15760 6480 16120 6540
rect 15800 6409 16120 6480
rect 14240 6100 15441 6380
rect 12300 5860 12360 6040
rect 12540 5860 12940 6040
rect 12300 5800 12600 5860
rect 12760 5600 12940 5860
rect 13800 6040 14100 6100
rect 13800 5860 13860 6040
rect 14040 6020 14100 6040
rect 14240 6020 14440 6100
rect 14040 5860 14440 6020
rect 13800 5800 14100 5860
rect 14260 5600 14440 5860
rect 15200 5980 15441 6100
rect -13100 5545 -12300 5600
rect -13100 3862 -13050 5545
rect -12860 5527 -12300 5545
rect -13100 3860 -13040 3862
rect -12860 3860 -12545 5527
rect -13100 3844 -12545 3860
rect -12355 3844 -12300 5527
rect -13100 3840 -12540 3844
rect -12360 3840 -12300 3844
rect -13100 3800 -12300 3840
rect -11600 5520 -11300 5600
rect -11600 3840 -11540 5520
rect -11360 3840 -11300 5520
rect -11600 3800 -11300 3840
rect -10600 5527 -10300 5600
rect -10600 3840 -10540 5527
rect -10350 3844 -10300 5527
rect -10360 3840 -10300 3844
rect -10600 3800 -10300 3840
rect -9600 5520 -9300 5600
rect -9600 3840 -9540 5520
rect -9360 3840 -9300 5520
rect -9600 3800 -9300 3840
rect -8600 5541 -7300 5600
rect -8600 5520 -8040 5541
rect -8600 3837 -8541 5520
rect -8351 3858 -8040 5520
rect -7850 5523 -7300 5541
rect -7850 3858 -7549 5523
rect -8351 3840 -7549 3858
rect -7359 3840 -7300 5523
rect -8351 3837 -7300 3840
rect -8600 3800 -7300 3837
rect -6900 5520 -6600 5600
rect -6900 3840 -6840 5520
rect -6660 3840 -6600 5520
rect -6900 3800 -6600 3840
rect -6200 5520 -5900 5600
rect -6200 3840 -6140 5520
rect -6200 3837 -6138 3840
rect -5948 3837 -5900 5520
rect -6200 3800 -5900 3837
rect -5500 5520 -5200 5600
rect -5500 3840 -5440 5520
rect -5260 3840 -5200 5520
rect -5500 3800 -5200 3840
rect -4800 5545 -3500 5600
rect -4800 5520 -4247 5545
rect -4800 3837 -4744 5520
rect -4554 3862 -4247 5520
rect -4057 5527 -3500 5545
rect -4057 3862 -3749 5527
rect -4554 3860 -4240 3862
rect -4060 3860 -3749 3862
rect -4554 3844 -3749 3860
rect -3559 3844 -3500 5527
rect -4554 3840 -3740 3844
rect -3560 3840 -3500 3844
rect -4554 3837 -3500 3840
rect -4800 3800 -3500 3837
rect -2300 5520 -2000 5600
rect -2300 3840 -2240 5520
rect -2060 3840 -2000 5520
rect -2300 3800 -2000 3840
rect -800 5520 -500 5600
rect -800 3840 -740 5520
rect -560 3840 -500 5520
rect -800 3800 -500 3840
rect 700 5541 2000 5600
rect 700 5523 1248 5541
rect 1438 5540 2000 5541
rect 700 3840 750 5523
rect 940 3858 1248 5523
rect 1440 5520 2000 5540
rect 1440 3860 1760 5520
rect 1438 3858 1760 3860
rect 940 3840 1760 3858
rect 700 3837 1763 3840
rect 1953 3837 2000 5520
rect 700 3800 2000 3837
rect 3200 5520 3500 5600
rect 3200 3840 3260 5520
rect 3440 3840 3500 5520
rect 3200 3800 3500 3840
rect 4700 5520 5000 5600
rect 4700 3840 4760 5520
rect 4940 3840 5000 5520
rect 4700 3800 5000 3840
rect 5200 5545 5500 5600
rect 5200 3862 5252 5545
rect 5442 3862 5500 5545
rect 5200 3860 5260 3862
rect 5440 3860 5500 3862
rect 5200 3800 5500 3860
rect 5700 5520 6000 5600
rect 5700 3840 5760 5520
rect 5940 3840 6000 5520
rect 5700 3800 6000 3840
rect 7200 5520 7500 5600
rect 7200 3840 7260 5520
rect 7440 3840 7500 5520
rect 7200 3800 7500 3840
rect 8700 5545 10000 5600
rect 8700 5527 9260 5545
rect 8700 3844 8755 5527
rect 8945 3860 9260 5527
rect 9450 5521 10000 5545
rect 9450 3862 9759 5521
rect 9440 3860 9759 3862
rect 8945 3844 9759 3860
rect 8700 3840 8760 3844
rect 8940 3843 9759 3844
rect 9942 3843 10000 5521
rect 8940 3840 9760 3843
rect 9940 3840 10000 3843
rect 8700 3800 10000 3840
rect 11200 5520 11500 5600
rect 11200 3840 11260 5520
rect 11440 3840 11500 5520
rect 11200 3800 11500 3840
rect 12700 5520 13000 5600
rect 12700 3840 12760 5520
rect 12940 3840 13000 5520
rect 12700 3800 13000 3840
rect 14200 5540 15000 5600
rect 14200 5520 14760 5540
rect 14940 5539 15000 5540
rect 14200 5518 14260 5520
rect 14200 3840 14253 5518
rect 14440 3860 14760 5520
rect 14944 3861 15000 5539
rect 15200 4840 15300 5980
rect 15831 5980 16081 6409
rect 16471 5973 16721 6338
rect 17111 5966 17361 6331
rect 17960 6400 18100 6760
rect 17960 6340 18001 6400
rect 18071 6340 18100 6400
rect 18300 6900 22700 6940
rect 18300 6760 20320 6900
rect 18300 6409 18420 6760
rect 19940 6409 20320 6760
rect 20720 6680 21080 6760
rect 20720 6620 20780 6680
rect 21020 6620 21080 6680
rect 20720 6560 21080 6620
rect 18300 6320 18321 6409
rect 18391 6320 18420 6409
rect 18711 5980 18961 6340
rect 19351 5980 19601 6209
rect 19465 5779 19601 5980
rect 19991 5980 20241 6409
rect 20311 6320 20320 6409
rect 20780 6320 21020 6560
rect 20631 5960 21100 6320
rect 20900 5740 21100 5960
rect 21260 5740 27720 5760
rect 20900 5300 27720 5740
rect 18640 4869 18709 4870
rect 15200 4440 15441 4840
rect 15760 4380 15761 4520
rect 15831 4379 16081 4820
rect 16360 4379 16401 4660
rect 16471 4379 16520 4660
rect 16791 4428 17041 4793
rect 17431 4441 17681 4806
rect 17480 4440 17640 4441
rect 17960 4379 18001 4600
rect 18071 4379 18120 4600
rect 15800 3960 16100 4379
rect 14940 3860 15000 3861
rect 14440 3840 15000 3860
rect 14200 3800 15000 3840
rect 15780 3880 16140 3960
rect 15780 3820 15840 3880
rect 16080 3820 16140 3880
rect 15780 3760 16140 3820
rect 16360 3680 16520 4379
rect 17960 4060 18120 4379
rect 18300 4379 18321 4620
rect 18391 4379 18420 4620
rect 18640 4380 18641 4869
rect 19031 4440 19281 4800
rect 19671 4440 19921 4800
rect 19991 4379 20241 4820
rect 20900 4820 21100 5300
rect 21260 5280 27720 5300
rect 20631 4460 21100 4820
rect 18300 4280 18420 4379
rect 19940 4280 20300 4379
rect 20540 4280 20900 4300
rect 18300 4220 20900 4280
rect 18300 4160 20600 4220
rect 20840 4160 20900 4220
rect 18300 4140 20900 4160
rect 20540 4100 20900 4140
rect 21520 4060 22120 4120
rect 17960 3860 21580 4060
rect 22060 3860 22120 4060
rect 21520 3820 22120 3860
rect 17420 3680 17740 3740
rect 16360 3480 17480 3680
rect 17680 3480 17740 3680
rect 17420 3440 17740 3480
<< viali >>
rect -13046 10340 -12860 10348
rect -13046 8663 -13040 10340
rect -13040 8663 -12860 10340
rect -12548 10340 -12362 10348
rect -12548 8663 -12540 10340
rect -12540 8663 -12362 10340
rect -11039 10340 -10853 10343
rect -11039 8660 -10860 10340
rect -10860 8660 -10853 10340
rect -10541 10340 -10355 10353
rect -10541 8668 -10540 10340
rect -10540 8668 -10360 10340
rect -10360 8668 -10355 10340
rect -10047 10340 -9861 10353
rect -10047 8668 -10040 10340
rect -10040 8668 -9861 10340
rect -11039 8658 -10853 8660
rect -6551 10340 -6365 10348
rect -6551 8663 -6540 10340
rect -6540 8663 -6365 10340
rect -2542 10340 -2356 10353
rect -2542 8668 -2540 10340
rect -2540 8668 -2360 10340
rect -2360 8668 -2356 10340
rect 1458 10340 1644 10348
rect 1458 8663 1460 10340
rect 1460 8663 1640 10340
rect 1640 8663 1644 10340
rect 4959 10340 5145 10353
rect 4959 8668 4960 10340
rect 4960 8668 5140 10340
rect 5140 8668 5145 10340
rect 6454 10340 6640 10343
rect 6454 8660 6460 10340
rect 6460 8660 6640 10340
rect 6957 10340 7143 10353
rect 6957 8668 6960 10340
rect 6960 8668 7140 10340
rect 7140 8668 7143 10340
rect 7460 10340 7646 10348
rect 7460 8663 7640 10340
rect 7640 8663 7646 10340
rect 6454 8658 6640 8660
rect 10458 10340 10644 10343
rect 10961 10340 11147 10343
rect 10458 8660 10460 10340
rect 10460 8660 10640 10340
rect 10640 8660 10644 10340
rect 10961 8660 11140 10340
rect 11140 8660 11147 10340
rect 11459 10340 11645 10353
rect 11459 8668 11460 10340
rect 11460 8668 11640 10340
rect 11640 8668 11645 10340
rect 10458 8658 10644 8660
rect 10961 8658 11147 8660
rect 14453 10340 14639 10353
rect 14956 10340 15142 10353
rect 14453 8668 14460 10340
rect 14460 8668 14639 10340
rect 14956 8668 14960 10340
rect 14960 8668 15140 10340
rect 15140 8668 15142 10340
rect 15459 10340 15645 10348
rect 15459 8663 15460 10340
rect 15460 8663 15640 10340
rect 15640 8663 15645 10340
rect 18457 10340 18643 10343
rect 18457 8660 18460 10340
rect 18460 8660 18640 10340
rect 18640 8660 18643 10340
rect 18951 10340 19137 10348
rect 19463 10340 19649 10348
rect 18951 8663 18960 10340
rect 18960 8663 19137 10340
rect 19463 8663 19640 10340
rect 19640 8663 19649 10340
rect 18457 8658 18643 8660
rect 20958 10340 21144 10348
rect 20958 8663 20960 10340
rect 20960 8663 21140 10340
rect 21140 8663 21144 10340
rect 4020 7242 4200 7442
rect 4020 6760 4200 6960
rect 6660 7240 6840 7440
rect 6660 6740 6840 6940
rect 10720 6742 10900 6942
rect 11720 7242 11900 7442
rect 23956 10340 24142 10348
rect 23956 8663 23960 10340
rect 23960 8663 24140 10340
rect 24140 8663 24142 10340
rect 24459 10340 24645 10353
rect 24459 8668 24460 10340
rect 24460 8668 24640 10340
rect 24640 8668 24645 10340
rect 24957 10340 25143 10353
rect 24957 8668 24960 10340
rect 24960 8668 25140 10340
rect 25140 8668 25143 10340
rect 26452 10340 26638 10348
rect 26955 10340 27141 10343
rect 26452 8663 26460 10340
rect 26460 8663 26638 10340
rect 26955 8660 26960 10340
rect 26960 8660 27140 10340
rect 27140 8660 27141 10340
rect 26955 8658 27141 8660
rect 15820 7620 16060 7780
rect 13440 7240 13620 7440
rect 21560 7240 22040 7440
rect 13440 6740 13620 6940
rect 15820 6540 16060 6600
rect -13050 5540 -12860 5545
rect -13050 3862 -13040 5540
rect -13040 3862 -12860 5540
rect -12545 5520 -12355 5527
rect -12545 3844 -12540 5520
rect -12540 3844 -12360 5520
rect -12360 3844 -12355 5520
rect -10540 5520 -10350 5527
rect -10540 3844 -10360 5520
rect -10360 3844 -10350 5520
rect -8040 5540 -7850 5541
rect -8541 3840 -8540 5520
rect -8540 3840 -8360 5520
rect -8360 3840 -8351 5520
rect -8040 3860 -7860 5540
rect -7860 3860 -7850 5540
rect -8040 3858 -7850 3860
rect -7549 5520 -7359 5523
rect -7549 3840 -7540 5520
rect -7540 3840 -7360 5520
rect -7360 3840 -7359 5520
rect -8541 3837 -8351 3840
rect -6138 3840 -5960 5520
rect -5960 3840 -5948 5520
rect -6138 3837 -5948 3840
rect -4247 5540 -4057 5545
rect -4744 3840 -4740 5520
rect -4740 3840 -4560 5520
rect -4560 3840 -4554 5520
rect -4247 3862 -4240 5540
rect -4240 3862 -4060 5540
rect -4060 3862 -4057 5540
rect -3749 5520 -3559 5527
rect -3749 3844 -3740 5520
rect -3740 3844 -3560 5520
rect -3560 3844 -3559 5520
rect -4744 3837 -4554 3840
rect 1248 5540 1438 5541
rect 750 5520 940 5523
rect 750 3840 760 5520
rect 760 3840 940 5520
rect 1248 3860 1260 5540
rect 1260 3860 1438 5540
rect 1248 3858 1438 3860
rect 1763 3840 1940 5520
rect 1940 3840 1953 5520
rect 1763 3837 1953 3840
rect 5252 5540 5442 5545
rect 5252 3862 5260 5540
rect 5260 3862 5440 5540
rect 5440 3862 5442 5540
rect 9260 5540 9450 5545
rect 8755 5520 8945 5527
rect 8755 3844 8760 5520
rect 8760 3844 8940 5520
rect 8940 3844 8945 5520
rect 9260 3862 9440 5540
rect 9440 3862 9450 5540
rect 9759 5520 9942 5521
rect 9759 3843 9760 5520
rect 9760 3843 9940 5520
rect 9940 3843 9942 5520
rect 14253 3840 14260 5518
rect 14260 3840 14436 5518
rect 14761 3861 14940 5539
rect 14940 3861 14944 5539
rect 17707 6003 17742 6355
rect 20780 6620 21020 6680
rect 15840 3820 16080 3880
rect 18658 4429 18697 4811
rect 20600 4160 20840 4220
rect 21580 3860 22060 4060
rect 17480 3480 17680 3680
<< metal1 >>
rect -13300 10353 27760 10400
rect -13300 10348 -10541 10353
rect -13300 8663 -13046 10348
rect -12860 8663 -12548 10348
rect -12362 10343 -10541 10348
rect -12362 8663 -11039 10343
rect -13300 8658 -11039 8663
rect -10853 8668 -10541 10343
rect -10355 8668 -10047 10353
rect -9861 10348 -2542 10353
rect -9861 8668 -6551 10348
rect -10853 8663 -6551 8668
rect -6365 8668 -2542 10348
rect -2356 10348 4959 10353
rect -2356 8668 1458 10348
rect -6365 8663 1458 8668
rect 1644 8668 4959 10348
rect 5145 10343 6957 10353
rect 5145 8668 6454 10343
rect 1644 8663 6454 8668
rect -10853 8658 6454 8663
rect 6640 8668 6957 10343
rect 7143 10348 11459 10353
rect 7143 8668 7460 10348
rect 6640 8663 7460 8668
rect 7646 10343 11459 10348
rect 7646 8663 10458 10343
rect 6640 8658 10458 8663
rect 10644 8658 10961 10343
rect 11147 8668 11459 10343
rect 11645 8668 14453 10353
rect 14639 8668 14956 10353
rect 15142 10348 24459 10353
rect 15142 8668 15459 10348
rect 11147 8663 15459 8668
rect 15645 10343 18951 10348
rect 15645 8663 18457 10343
rect 11147 8658 18457 8663
rect 18643 8663 18951 10343
rect 19137 8663 19463 10348
rect 19649 8663 20958 10348
rect 21144 8663 23956 10348
rect 24142 8668 24459 10348
rect 24645 8668 24957 10353
rect 25143 10348 27760 10353
rect 25143 8668 26452 10348
rect 24142 8663 26452 8668
rect 26638 10343 27760 10348
rect 26638 8663 26955 10343
rect 18643 8658 26955 8663
rect 27141 8658 27760 10343
rect -13300 8640 27760 8658
rect -13300 8600 27400 8640
rect 14600 8000 17000 8220
rect 3960 7460 4260 7502
rect 6600 7460 6900 7500
rect 3960 7442 6900 7460
rect 3960 7242 4020 7442
rect 4200 7440 6900 7442
rect 4200 7260 6660 7440
rect 4200 7242 4260 7260
rect 3960 7202 4260 7242
rect 6600 7240 6660 7260
rect 6840 7240 6900 7440
rect 6600 7200 6900 7240
rect 11660 7460 11960 7502
rect 13380 7460 13680 7500
rect 11660 7442 13680 7460
rect 11660 7242 11720 7442
rect 11900 7440 13680 7442
rect 11900 7260 13440 7440
rect 11900 7242 11960 7260
rect 11660 7202 11960 7242
rect 13380 7240 13440 7260
rect 13620 7240 13680 7440
rect 13380 7200 13680 7240
rect 3960 6960 4260 7020
rect 6600 6960 6900 7000
rect 3960 6760 4020 6960
rect 4200 6940 6900 6960
rect 4200 6760 6660 6940
rect 3960 6720 4260 6760
rect 6600 6740 6660 6760
rect 6840 6740 6900 6940
rect 6600 6700 6900 6740
rect 10660 6960 10960 7002
rect 13380 6960 13680 7000
rect 10660 6942 13680 6960
rect 10660 6742 10720 6942
rect 10900 6940 13680 6942
rect 10900 6760 13440 6940
rect 10900 6742 10960 6760
rect 10660 6702 10960 6742
rect 13380 6740 13440 6760
rect 13620 6740 13680 6940
rect 13380 6700 13680 6740
rect 14600 5600 15060 8000
rect 15760 7780 16120 7860
rect 15760 7620 15820 7780
rect 16060 7620 16120 7780
rect 15760 7540 16120 7620
rect 15840 6680 16040 7540
rect 16660 7320 17000 8000
rect 21500 7440 22100 7500
rect 16660 7100 21020 7320
rect 21500 7240 21560 7440
rect 22040 7240 22100 7440
rect 21500 7200 22100 7240
rect 20760 6760 21020 7100
rect 20720 6680 21080 6760
rect 15760 6600 16120 6680
rect 18526 6672 18579 6673
rect 15760 6540 15820 6600
rect 16060 6540 16120 6600
rect 15760 6480 16120 6540
rect 17674 6588 18579 6672
rect 17674 6393 17768 6588
rect 17681 6355 17751 6393
rect 17681 6003 17707 6355
rect 17742 6003 17751 6355
rect 17681 5922 17751 6003
rect -13300 5545 15100 5600
rect -13300 3862 -13050 5545
rect -12860 5541 -4247 5545
rect -12860 5527 -8040 5541
rect -12860 3862 -12545 5527
rect -13300 3844 -12545 3862
rect -12355 3844 -10540 5527
rect -10350 5520 -8040 5527
rect -10350 3844 -8541 5520
rect -13300 3837 -8541 3844
rect -8351 3858 -8040 5520
rect -7850 5523 -4247 5541
rect -7850 3858 -7549 5523
rect -8351 3840 -7549 3858
rect -7359 5520 -4247 5523
rect -7359 3840 -6138 5520
rect -8351 3837 -6138 3840
rect -5948 3837 -4744 5520
rect -4554 3862 -4247 5520
rect -4057 5541 5252 5545
rect -4057 5527 1248 5541
rect -4057 3862 -3749 5527
rect -4554 3844 -3749 3862
rect -3559 5523 1248 5527
rect -3559 3844 750 5523
rect -4554 3840 750 3844
rect 940 3858 1248 5523
rect 1438 5520 5252 5541
rect 1438 3858 1763 5520
rect 940 3840 1763 3858
rect -4554 3837 1763 3840
rect 1953 3862 5252 5520
rect 5442 5527 9260 5545
rect 5442 3862 8755 5527
rect 1953 3844 8755 3862
rect 8945 3862 9260 5527
rect 9450 5539 15100 5545
rect 9450 5521 14761 5539
rect 9450 3862 9759 5521
rect 8945 3844 9759 3862
rect 1953 3843 9759 3844
rect 9942 5518 14761 5521
rect 9942 3843 14253 5518
rect 1953 3840 14253 3843
rect 14436 3861 14761 5518
rect 14944 3861 15100 5539
rect 18510 4832 18579 6588
rect 20720 6620 20780 6680
rect 21020 6620 21080 6680
rect 20720 6560 21080 6620
rect 21600 6420 22020 7200
rect 22920 5880 27160 6420
rect 21560 5820 22060 5860
rect 21520 5180 22000 5200
rect 24000 5180 26080 5880
rect 21520 5160 26080 5180
rect 18640 4832 18709 4870
rect 18510 4811 18709 4832
rect 18510 4429 18658 4811
rect 18697 4429 18709 4811
rect 18510 4380 18709 4429
rect 21520 4660 26100 5160
rect 21520 4640 25860 4660
rect 18510 4379 18707 4380
rect 20540 4220 20900 4300
rect 20540 4160 20600 4220
rect 20840 4160 20900 4220
rect 20540 4100 20900 4160
rect 14436 3840 15100 3861
rect 1953 3837 15100 3840
rect -13300 3800 15100 3837
rect 15780 3900 16140 3960
rect 20600 3900 20900 4100
rect 15780 3880 20900 3900
rect 15780 3820 15840 3880
rect 16080 3820 20900 3880
rect 21520 4060 22240 4640
rect 21520 3860 21580 4060
rect 22060 4000 22240 4060
rect 22060 3860 22120 4000
rect 21520 3820 22120 3860
rect 15780 3800 20900 3820
rect 15780 3760 16140 3800
rect 17420 3680 17740 3740
rect 26780 3680 27400 4880
rect 17420 3480 17480 3680
rect 17680 3500 27400 3680
rect 17680 3480 17740 3500
rect 17420 3440 17740 3480
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 1 1288
timestamp 1665323087
transform 1 0 21244 0 1 4202
box 0 0 1340 1340
<< labels >>
flabel poly -9700 8100 -9700 8100 0 FreeSans 1600 0 0 0 MSU
flabel poly 9300 8100 9300 8100 0 FreeSans 1600 0 0 0 a
flabel poly -6500 6580 -6500 6580 0 FreeSans 1600 0 0 0 b
flabel locali 11220 7460 11220 7460 0 FreeSans 1600 0 0 0 VD1
flabel locali 7420 6960 7420 6960 0 FreeSans 1600 0 0 0 VDR
flabel locali 21180 3960 21180 3960 0 FreeSans 1600 0 0 0 VD2
flabel metal1 18380 3580 18380 3580 0 FreeSans 1600 0 0 0 VD3
flabel locali 27760 7700 27760 7700 0 FreeSans 1600 0 0 0 Vref
rlabel metal1 -13300 9500 -13300 9500 7 VDD
rlabel metal1 -13300 4700 -13300 4700 7 GND
<< end >>
